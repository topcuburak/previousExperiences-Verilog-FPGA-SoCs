library verilog;
use verilog.vl_types.all;
entity hw_2_vlg_vec_tst is
end hw_2_vlg_vec_tst;
