library verilog;
use verilog.vl_types.all;
entity hw_2_vlg_check_tst is
    port(
        out_1           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hw_2_vlg_check_tst;
